module Instruction_Memory
(
	input [63:0] Inst_Address,
	output reg [31:0] Instruction
);
	reg [7:0] inst_mem [147:0];
	
initial
	begin
		inst_mem[0]  = 8'h93; // more explanation of code in part 1
		inst_mem[1]  = 8'h05;
		inst_mem[2]  = 8'h60;
		inst_mem[3]  = 8'h00;
		inst_mem[4]  = 8'h93;
		inst_mem[5]  = 8'h0E;
		inst_mem[6]  = 8'h60;
		inst_mem[7]  = 8'h00;
		inst_mem[8]  = 8'h13;
		inst_mem[9]  = 8'h0F;
		inst_mem[10] = 8'h00;
		inst_mem[11] = 8'h00;
		inst_mem[12] = 8'h13;
		inst_mem[13] = 8'h0F;
		inst_mem[14] = 8'h00;
		inst_mem[15] = 8'h00;
		inst_mem[16] = 8'h13;
		inst_mem[17] = 8'h0E;
		inst_mem[18] = 8'h60;
		inst_mem[19] = 8'h00;
		inst_mem[20] = 8'h23;
		inst_mem[21] = 8'h20;
		inst_mem[22] = 8'hBF;
		inst_mem[23] = 8'h10;
		inst_mem[24] = 8'h93;
		inst_mem[25] = 8'h8F;
		inst_mem[26] = 8'h1F;
		inst_mem[27] = 8'h00;
		inst_mem[28] = 8'h13;
		inst_mem[29] = 8'h0F;
		inst_mem[30] = 8'h8F;
		inst_mem[31] = 8'h00;
		inst_mem[32] = 8'h93;
		inst_mem[33] = 8'h85;
		inst_mem[34] = 8'hF5;
		inst_mem[35] = 8'hFF;
		inst_mem[36] = 8'h63;
		inst_mem[37] = 8'h04;
		inst_mem[38] = 8'hFE;
		inst_mem[39] = 8'h01;
		inst_mem[40] = 8'hE3;
		inst_mem[41] = 8'h06;
		inst_mem[42] = 8'h00;
		inst_mem[43] = 8'hFE;
		inst_mem[44] = 8'h13;
		inst_mem[45] = 8'h0F;
		inst_mem[46] = 8'h00;
		inst_mem[47] = 8'h00;
		inst_mem[48] = 8'h93;
		inst_mem[49] = 8'h0F;
		inst_mem[50] = 8'h0F;
		inst_mem[51] = 8'h00;
		inst_mem[52] = 8'h93;
		inst_mem[53] = 8'h0E;
		inst_mem[54] = 8'h00;
		inst_mem[55] = 8'h00;
		inst_mem[56] = 8'h93;
		inst_mem[57] = 8'h05;
		inst_mem[58] = 8'h60;
		inst_mem[59] = 8'h00;
		inst_mem[60] = 8'h63;
		inst_mem[61] = 8'h8C;
		inst_mem[62] = 8'hE5;
		inst_mem[63] = 8'h05;
		inst_mem[64] = 8'h33;
		inst_mem[65] = 8'h85;
		inst_mem[66] = 8'h0E;
		inst_mem[67] = 8'h00;
		inst_mem[68] = 8'h93;
		inst_mem[69] = 8'h0F;
		inst_mem[70] = 8'h1F;
		inst_mem[71] = 8'h00;
		inst_mem[72] = 8'h13;
		inst_mem[73] = 8'h8E;
		inst_mem[74] = 8'h8E;
		inst_mem[75] = 8'h00;
		inst_mem[76] = 8'h63;
		inst_mem[77] = 8'h88;
		inst_mem[78] = 8'hBF;
		inst_mem[79] = 8'h02;
		inst_mem[80] = 8'h83;
		inst_mem[81] = 8'h27;
		inst_mem[82] = 8'h0E;
		inst_mem[83] = 8'h10;
		inst_mem[84] = 8'h03;
		inst_mem[85] = 8'h28;
		inst_mem[86] = 8'h05;
		inst_mem[87] = 8'h10;
		inst_mem[88] = 8'h63;
		inst_mem[89] = 8'hCE;
		inst_mem[90] = 8'h07;
		inst_mem[91] = 8'h01;
		inst_mem[92] = 8'h93;
		inst_mem[93] = 8'h8F;
		inst_mem[94] = 8'h1F;
		inst_mem[95] = 8'h00;
		inst_mem[96] = 8'h13;
		inst_mem[97] = 8'h0E;
		inst_mem[98] = 8'h8E;
		inst_mem[99] = 8'h00;
		inst_mem[100] = 8'hE3;
		inst_mem[101] = 8'h04;
		inst_mem[102] = 8'h00;
		inst_mem[103] = 8'hFC;
		inst_mem[104] = 8'h13;
		inst_mem[105] = 8'h0F;
		inst_mem[106] = 8'h1F;
		inst_mem[107] = 8'h00;
		inst_mem[108] = 8'h13;
		inst_mem[109] = 8'h0E;
		inst_mem[110] = 8'h8E;
		inst_mem[111] = 8'h00;
		inst_mem[112] = 8'hE3;
		inst_mem[113] = 8'h06;
		inst_mem[114] = 8'h00;
		inst_mem[115] = 8'hFC;
		inst_mem[116] = 8'h13;
		inst_mem[117] = 8'h05;
		inst_mem[118] = 8'h0E;
		inst_mem[119] = 8'h00;
		inst_mem[120] = 8'hE3;
		inst_mem[121] = 8'h02;
		inst_mem[122] = 8'h00;
		inst_mem[123] = 8'hFE;
		inst_mem[124] = 8'h83;
		inst_mem[125] = 8'h26;
		inst_mem[126] = 8'h05;
		inst_mem[127] = 8'h10;
		inst_mem[128] = 8'h03;
		inst_mem[129] = 8'hA7;
		inst_mem[130] = 8'h0E;
		inst_mem[131] = 8'h10;
		inst_mem[132] = 8'h23;
		inst_mem[133] = 8'hA0;
		inst_mem[134] = 8'hDE;
		inst_mem[135] = 8'h10;
		inst_mem[136] = 8'h23;
		inst_mem[137] = 8'h20;
		inst_mem[138] = 8'hE5;
		inst_mem[139] = 8'h10;
		inst_mem[140] = 8'h93;
		inst_mem[141] = 8'h8E;
		inst_mem[142] = 8'h8E;
		inst_mem[143] = 8'h00;
		inst_mem[144] = 8'hE3;
		inst_mem[145] = 8'h06;
		inst_mem[146] = 8'h00;
		inst_mem[147] = 8'hFC;
	end
	
	always @(Inst_Address)
	begin
		Instruction={inst_mem[Inst_Address+3],inst_mem[Inst_Address+2],inst_mem[Inst_Address+1],inst_mem[Inst_Address]};
	end
endmodule
