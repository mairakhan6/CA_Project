module EX_MEM(
    input clk,                     // Clock signal
    input Flush,                   // Flush control signal
    input RegWrite,                // Control signal for enabling register write
    input MemtoReg,                // Control signal for selecting memory or ALU result for register write
    input Branch,                  // Control signal for branch instruction
    input Zero,                    // Control signal indicating the ALU result is zero
    input MemWrite,                // Control signal for memory write
    input MemRead,                 // Control signal for memory read
    input is_greater,              // Control signal indicating the comparison result of the ALU operation
    input [63:0] immvalue_added_pc, // Immediate value added to the program counter
    input [63:0] ALU_result,       // Result of the ALU operation
    input [63:0] WriteData,        // Data to be written to memory or register file
    input [3:0] function_code,     // Function code for ALU operation
    input [4:0] destination_reg,   // Destination register for register write

    output reg RegWrite_out,       // Output signal for enabling register write
    output reg MemtoReg_out,       // Output signal for selecting memory or ALU result for register write
    output reg Branch_out,         // Output signal for branch instruction
    output reg Zero_out,           // Output signal indicating the ALU result is zero
    output reg MemWrite_out,       // Output signal for memory write
    output reg MemRead_out,        // Output signal for memory read
    output reg is_greater_out,     // Output signal indicating the comparison result of the ALU operation
    output reg [63:0] immvalue_added_pc_out, // Output signal for immediate value added to the program counter
    output reg [63:0] ALU_result_out,       // Output signal for the ALU result
    output reg [63:0] WriteData_out,        // Output signal for data to be written to memory or register file
    output reg [3:0] function_code_out,     // Output signal for function code for ALU operation
    output reg [4:0] destination_reg_out    // Output signal for destination register for register write
);

    // Assign output values based on control signals
    always @(posedge clk) begin
        if (Flush) begin
            // Reset output values when flush signal is active
            RegWrite_out = 0;
            MemtoReg_out = 0;
            Branch_out = 0;
            Zero_out = 0;
            is_greater_out = 0;
            MemWrite_out = 0;
            MemRead_out = 0;
            immvalue_added_pc_out = 0;
            ALU_result_out = 0;
            WriteData_out = 0;
            function_code_out = 0;
            destination_reg_out = 0;
        end 
        else begin
            // Assign output values based on input signals
            RegWrite_out = RegWrite;
            MemtoReg_out = MemtoReg;
            Branch_out = Branch;
            Zero_out = Zero;
            is_greater_out = is_greater;
            MemWrite_out = MemWrite;
            MemRead_out = MemRead;
            immvalue_added_pc_out = immvalue_added_pc;
            ALU_result_out = ALU_result;
            WriteData_out = WriteData;
            function_code_out = function_code;
            destination_reg_out = destination_reg;
        end
    end

endmodule